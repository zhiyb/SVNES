`include "config.h"

module cpu (
);

endmodule
