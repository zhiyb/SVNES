`include "config.h"

module pc (
);

endmodule
